resp_tx.vhd